/***************************************
#
#			Filename:decoder.sv
#
#			Developer:ske
#			Description:---
#			CreatTime:2021-09-27 22:22:20
#
***************************************/
module decoder(
    input logic clk_i,
    input logic rst_ni,
    // from IF-ID pipeline register
    input logic [31:0] instr_rdata_i, //指令数据输入，来自指令ram
    // immediates
    //output logic 
    // register file
    output logic 
);


endmodule

