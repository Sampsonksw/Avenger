/***************************************
#
#			Filename:milano.sv
#
#			Developer:ske
#			Description:---
#			CreatTime:2021-09-29 15:09:11
#
***************************************/

module milano(
        input  logic clk_i,
        input  logic rst_ni,
        //input from boot sel
        input  logic [31:0] boot_addr_i,
        //output to system bus
        output logic [31:0] instr_addr_o
);




/********** if stage unit  ***********/


/********** id stage unit  **********/

/********** ex stage unit  **********/

endmodule
